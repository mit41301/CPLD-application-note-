library verilog;
use verilog.vl_types.all;
entity SPI_to_I2C_test is
end SPI_to_I2C_test;
