library verilog;
use verilog.vl_types.all;
entity SPI_master_test is
end SPI_master_test;
