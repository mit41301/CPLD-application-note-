library verilog;
use verilog.vl_types.all;
entity test_ufm_memory is
end test_ufm_memory;
